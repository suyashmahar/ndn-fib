// `ifndef _my_incl_vh_
//  `define _my_incl_vh_
// 
//  `define NULL 0
// 
//  // Defines global Parameters
//  `define WORD_SIZE = 64;
//  `define POINTER_SIZE = 16;
//  `define MAX_NAME_LENGTH = 16; // max length of name in words
// `endif
